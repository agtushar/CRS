../globals.vhd